library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

use work.constants.ALL;

entity VGA is
	port (
		clk_i : in STD_LOGIC;
		rst_ni : in STD_LOGIC;

		hsync_o : out STD_LOGIC;
		vsync_o : out STD_LOGIC;

		registers_i : in reg_t;
		registers_fp_i : in reg_t;

		fcsr_i : in STD_LOGIC_VECTOR (7 downto 0);

		pc_i : in STD_LOGIC_VECTOR (63 downto 0);
		rgb_o : out STD_LOGIC_VECTOR (11 downto 0));
end VGA;

architecture behavioral of VGA is
    
    constant HSP : integer := 96; 
    constant TH : integer := 800;
    constant HDT : integer := 640;
    constant HBP : integer := 48;
    constant HFP : integer := 16;

    constant VSP : integer := 2; 
    constant TV : integer := 521;
    constant VDT : integer := 480;
    constant VBP : integer := 29;
    constant VFP : integer := 10;

    type char_ram is array (0 to 79) of STD_LOGIC_VECTOR (639 downto 0);    
    signal frame_buffer : char_ram := (
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2C2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2D",
        X"2B2929292929292929292929292929291113170E100E16292929292929292929292929292929292B292929292929292929292929290F12140A171113102915141113172929292929292929292929292B",
        X"2B2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2B",
        X"2B291319201C2929291326201A1C232929292929292929292918191F261C2929292929292929292B291319201C292929291326201A1C232929292929292929292918191F261C2929292929292929292B",
        X"2B2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2B",
        X"2B29281C23212929292929002929292929292900270000000000000000000000000000000029292B291D250029292929292929002929292929292900270000000000000000000000000000000029292B",
        X"2B29231929292929292929012929292929292900270000000000000000000000000000000029292B291D250129292929292929012929292929292900270000000000000000000000000000000029292B",
        X"2B29242229292929292929022929292929292900270000000000000000000000000000000029292B291D250229292929292929022929292929292900270000000000000000000000000000000029292B",
        X"2B291E2229292929292929032929292929292900270000000000000000000000000000000029292B291D250329292929292929032929292929292900270000000000000000000000000000000029292B",
        X"2B29252229292929292929042929292929292900270000000000000000000000000000000029292B291D250429292929292929042929292929292900270000000000000000000000000000000029292B",
        X"2B29250029292929292929052929292929292900270000000000000000000000000000000029292B291D250529292929292929052929292929292900270000000000000000000000000000000029292B",
        X"2B29250129292929292929062929292929292900270000000000000000000000000000000029292B291D250629292929292929062929292929292900270000000000000000000000000000000029292B",
        X"2B29250229292929292929072929292929292900270000000000000000000000000000000029292B291D250729292929292929072929292929292900270000000000000000000000000000000029292B",
        X"2B29240029292929292929082929292929292900270000000000000000000000000000000029292B291D240029292929292929082929292929292900270000000000000000000000000000000029292B",
        X"2B29240129292929292929092929292929292900270000000000000000000000000000000029292B291D240129292929292929092929292929292900270000000000000000000000000000000029292B",
        X"2B29190029292929292929010029292929292900270000000000000000000000000000000029292B291D190029292929292929010029292929292900270000000000000000000000000000000029292B",
        X"2B29190129292929292929010129292929292900270000000000000000000000000000000029292B291D190129292929292929010129292929292900270000000000000000000000000000000029292B",
        X"2B29190229292929292929010229292929292900270000000000000000000000000000000029292B291D190229292929292929010229292929292900270000000000000000000000000000000029292B",
        X"2B29190329292929292929010329292929292900270000000000000000000000000000000029292B291D190329292929292929010329292929292900270000000000000000000000000000000029292B",
        X"2B29190429292929292929010429292929292900270000000000000000000000000000000029292B291D190429292929292929010429292929292900270000000000000000000000000000000029292B",
        X"2B29190529292929292929010529292929292900270000000000000000000000000000000029292B291D190529292929292929010529292929292900270000000000000000000000000000000029292B",
        X"2B29190629292929292929010629292929292900270000000000000000000000000000000029292B291D190629292929292929010629292929292900270000000000000000000000000000000029292B",
        X"2B29190729292929292929010729292929292900270000000000000000000000000000000029292B291D190729292929292929010729292929292900270000000000000000000000000000000029292B",
        X"2B29240229292929292929010829292929292900270000000000000000000000000000000029292B291D240229292929292929010829292929292900270000000000000000000000000000000029292B",
        X"2B29240329292929292929010929292929292900270000000000000000000000000000000029292B291D240329292929292929010929292929292900270000000000000000000000000000000029292B",
        X"2B29240429292929292929020029292929292900270000000000000000000000000000000029292B291D240429292929292929020029292929292900270000000000000000000000000000000029292B",
        X"2B29240529292929292929020129292929292900270000000000000000000000000000000029292B291D240529292929292929020129292929292900270000000000000000000000000000000029292B",
        X"2B29240629292929292929020229292929292900270000000000000000000000000000000029292B291D240629292929292929020229292929292900270000000000000000000000000000000029292B",
        X"2B29240729292929292929020329292929292900270000000000000000000000000000000029292B291D240729292929292929020329292929292900270000000000000000000000000000000029292B",
        X"2B29240829292929292929020429292929292900270000000000000000000000000000000029292B291D240829292929292929020429292929292900270000000000000000000000000000000029292B",
        X"2B29240929292929292929020529292929292900270000000000000000000000000000000029292B291D240929292929292929020529292929292900270000000000000000000000000000000029292B",
        X"2B29240100292929292929020629292929292900270000000000000000000000000000000029292B291D240100292929292929020629292929292900270000000000000000000000000000000029292B",
        X"2B29240101292929292929020729292929292900270000000000000000000000000000000029292B291D240101292929292929020729292929292900270000000000000000000000000000000029292B",
        X"2B29250329292929292929020829292929292900270000000000000000000000000000000029292B291D250829292929292929020829292929292900270000000000000000000000000000000029292B",
        X"2B29250429292929292929020929292929292900270000000000000000000000000000000029292B291D250929292929292929020929292929292900270000000000000000000000000000000029292B",
        X"2B29250529292929292929030029292929292900270000000000000000000000000000000029292B291D250100292929292929030029292929292900270000000000000000000000000000000029292B",
        X"2B29250629292929292929030129292929292900270000000000000000000000000000000029292B291D250101292929292929030129292929292900270000000000000000000000000000000029292B",
        X"2B2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2B2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2B",
        X"2B29150C29292929292929292929292929292900270000000000000000000000000000000029292B291D1B2423292929292929292929292929292929292929002700000000000000002929292929292B",
        X"2E2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2F",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929",
        X"2929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929292929"
    );
    
    function to_oct(reg : STD_LOGIC_VECTOR) return STD_LOGIC_VECTOR is
        variable oct : STD_LOGIC_VECTOR (2 * reg'length - 1 downto 0);
    begin
        for i in 0 to reg'length/4 - 1 loop
            oct(i * 8 + 7 downto i * 8) := X"0" & reg(i * 4 + 3 downto i * 4);
        end loop;
        return oct;
    end function;
    
	
    signal pixel_clk, hsync_reg, vsync_reg, display : STD_LOGIC := '0';
    signal counter : STD_LOGIC_VECTOR (1 downto 0) := "00";
 
    signal hcount, vcount : STD_LOGIC_VECTOR (9 downto 0) := (others => '0');       
 
    signal row_font : STD_LOGIC_VECTOR (10 downto 0);
    signal row, column : STD_LOGIC_VECTOR (9 downto 0);

    signal font_data : STD_LOGIC_VECTOR (7 downto 0);
 
    component font_ROM is
        port ( row_i : in STD_LOGIC_VECTOR (10 downto 0);
               data_o : out STD_LOGIC_VECTOR (7 downto 0));
    end component font_ROM;
 
begin

	PRESCALER : process (clk_i)
	begin
		if rising_edge(clk_i) then
			if rst_ni = '0' then
				counter <= "00";
				pixel_clk <= '0';
				else
				if counter = 3 then
					counter <= "00";
					pixel_clk <= '1';
				else
					counter <= counter + 1;
					pixel_clk <= '0';
				end if;
			end if;
		end if;
	end process;

	COUNTERS : process (clk_i)
	begin
		if rising_edge(clk_i) then
			if rst_ni = '0' then
				hcount <= (others => '0');
				vcount <= (others => '0');
				else
				if pixel_clk = '1' then
					if hcount = TH - 1 then
						hcount <= (others => '0');
						if vcount = TV - 1 then
							vcount <= (others => '0');
						else
							vcount <= vcount + 1;
						end if;
					else
						hcount <= hcount + 1;
					end if;
				end if;
			end if;
		end if;
	end process;

	HSYNC : process (clk_i)
	begin
		if rising_edge(clk_i) then
			if hcount < HDT + HFP or hcount >= HDT + HFP + HSP then
 				hsync_reg <= '1';
			else
				hsync_reg <= '0';
			end if;
		end if;
	end process;

	VSYNC : process (clk_i)
	begin
		if rising_edge(clk_i) then
			if vcount < VDT + VFP or vcount >= VDT + VFP + VSP then
				vsync_reg <= '1';
				else
				vsync_reg <= '0';
			end if;
		end if;
	end process;

	row <= vcount when vcount < VDT else (others => '0');
	column <= hcount when hcount < HDT else (others => '0');
	display <= '1' when hcount < HDT and vcount < VDT else '0';

	DISPLAY_REGISTERS_CONTENTS : for i in 0 to 31 generate
		frame_buffer(i + 25)(471 downto 344) <= to_oct(registers_i(i));
		frame_buffer(i + 25)(151 downto 24) <= to_oct(registers_fp_i(i));
	end generate;

	frame_buffer(58)(471 downto 344) <= to_oct(pc_i);
	frame_buffer(58)(71 downto 56) <= to_oct(fcsr_i);

	hsync_o <= hsync_reg;
	vsync_o <= vsync_reg;

	row_font <= frame_buffer(conv_integer(row(8 downto 3)))(639 - 8 * conv_integer(column(9 downto 3)) downto 632 - 8 * conv_integer(column(9 downto 3))) & row(2 downto 0);

	rgb_o <= (others => '1') when font_data(7 - conv_integer(column(2 downto 0))) = '1' and display = '1' else (others => '0');

	FONT : font_ROM
	port map(
		row_i => row_font,
		data_o => font_data
	);
   
end behavioral;