-- https://github.com/martimdfneves/ECT/blob/ba39a5b4e36656bcb0fa5b26c46a69df45b93914/1%20ano/2%20semestre/LSD/lsd_support/vhdl_code/font_8x8_bold.vhd

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity font_ROM is
    port ( 
		row_i : in STD_LOGIC_VECTOR (10 downto 0);
        data_o : out STD_LOGIC_VECTOR (7 downto 0));
end font_ROM;

architecture behavioral of font_ROM is
    type rom_type is array (0 to 383) of STD_LOGIC_VECTOR (7 downto 0);
    signal rom : rom_type := (
        -- 0 0x00
        "01111100",
        "11000110",
        "11000110", 
        "11000110",
        "11000110",
        "11000110",
        "01111100",
        --1
        "00000000",
        "00110000",
        "01110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "11111100",
        "00000000",
        --2
        "01111000",
        "11001100",
        "00001100",
        "00111000",
        "01100000",
        "11001100",
        "11111100",
        "00000000",
        --3
        "01111000",
        "11001100",
        "00001100",
        "00111000",
        "00001100",
        "11001100",
        "01111000",
        "00000000",
        --4
        "00011100",
        "00111100",
        "01101100",
        "11001100",
        "11111110",
        "00001100",
        "00011110",
        "00000000",
        --5
        "11111100",
        "11000000",
        "11111000",
        "00001100",
        "00001100",
        "11001100",
        "01111000",
        "00000000",
        --6
        "00111000",
        "01100000",
        "11000000",
        "11111000",
        "11001100",
        "11001100",
        "01111000",
        "00000000",
        --7
        "11111100",
        "11001100",
        "00001100",
        "00011000",
        "00110000",
        "00110000",
        "00110000",
        "00000000",
        --8
        "01111000",
        "11001100",
        "11001100",
        "01111000",
        "11001100",
        "11001100",
        "01111000",
        "00000000",
        --9
        "01111000",
        "11001100",
        "11001100",
        "01111100",
        "00001100",
        "00011000",
        "01110000",
        "00000000",
        --A
        "00110000",
        "01111000",
        "11001100",
        "11001100",
        "11111100",
        "11001100",
        "11001100",
        "00000000",
        --B
        "11111100",
        "01100110",
        "01100110",
        "01111100",
        "01100110",
        "01100110",
        "11111100",
        "00000000",
        --C
        "00111100",
        "01100110",
        "11000000",
        "11000000",
        "11000000",
        "01100110",
        "00111100",
        "00000000",
        --D
        "11111000",
        "01101100",
        "01100110",
        "01100110",
        "01100110",
        "01101100",
        "11111000",
        "00000000",
        --E
        "11111110",
        "01100010",
        "01101000",
        "01111000",
        "01101000",
        "01100010",
        "11111110",
        "00000000",
        --F
        "11111110",
        "01100010",
        "01101000",
        "01111000",
        "01101000",
        "01100000",
        "11110000",
        "00000000", 
       --[0x10] G
        "00111100",
        "01100110",
        "11000000",
        "11000000",
        "11001110",
        "01100110",
        "00111110",
        "00000000",
       -- [0x11] I
        "01111000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "01111000",
        "00000000",
      -- [0x12] L
        "11110000",
        "01100000",
        "01100000",
        "01100000",
        "01100010",
        "01100110",
        "11111110",
        "00000000",   
        -- [ 0x13] N
        "11000110",
        "11100110",
        "11110110",
        "11011110",
        "11001110",
        "11000110",
        "11000110",
        "00000000",
      -- [0x14] O
        "00111000",
        "01101100",
        "11000110",
        "11000110",
        "11000110",
        "01101100",
        "00111000",
        "00000000",
      -- [0X15] P
        "11111100",
        "01100110",
        "01100110",
        "01111100",
        "01100000",
        "01100000",
        "11110000",
        "00000000",
      -- [0x16] R
        "11111100",
        "01100110",
        "01100110",
        "01111100",
        "01101100",
        "01100110",
        "11100110",
        "00000000",
      -- [0x17] T
        "11111100",
        "10110100",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "01111000",
        "00000000", 
       -- [ 0x18] V
        "11001100",
        "11001100",
        "11001100",
        "11001100",
        "11001100",
        "01111000",
        "00110000",
        "00000000",
     -- [ 0x19] a
        "00000000",
        "00000000",
        "01111000",
        "00001100",
        "01111100",
        "11001100",
        "01110110",
        "00000000",
     -- [ 0x1A] b
        "11100000",
        "01100000",
        "01100000",
        "01111100",
        "01100110",
        "01100110",
        "11011100",
        "00000000",
    -- [ 0x1B] c   
        "00000000",
        "00000000",
        "01111000",
        "11001100",
        "11000000",
        "11001100",
        "01111000",
        "00000000",
      -- [0x1C] e
        "00000000",
        "00000000",
        "01111000",
        "11001100",
        "11111100",
        "11000000",
        "01111000",
        "00000000",
     -- [0x1D] f
        "00111000",
        "01101100",
        "01100000",
        "11110000",
        "01100000",
        "01100000",
        "11110000",
        "00000000",
       -- [0x1E] g
        "00000000",
        "00000000",
        "01110110",
        "11001100",
        "11001100",
        "01111100",
        "00001100",
        "11111000",
      -- [0x1F] l
        "01110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "01111000",
        "00000000",
       -- [0x20] m
        "00000000",
        "00000000",
        "11001100",
        "11111110",
        "11111110",
        "11010110",
        "11000110",
        "00000000",
        -- [0x21] o
        "00000000",
        "00000000",
        "01111000",
        "11001100",
        "11001100",
        "11001100",
        "01111000",
        "00000000",
       -- [0x22] p
        "00000000",
        "00000000",
        "11011100",
        "01100110",
        "01100110",
        "01111100",
        "01100000",
        "11110000",
       -- [0x23] r
        "00000000",
        "00000000",
        "11011100",
        "01110110",
        "01100110",
        "01100000",
        "11110000",
        "00000000",
       -- [0x24] s
        "00000000",
        "00000000",
        "01111100",
        "11000000",
        "01111000",
        "00001100",
        "11111000",
        "00000000",
       -- [0x25] t
        "00010000",
        "00110000",
        "01111100",
        "00110000",
        "00110000",
        "00110100",
        "00011000",
        "00000000",
       -- [0x26] u
        "00000000",
        "00000000",
        "11001100",
        "11001100",
        "11001100",
        "11001100",
        "01110110",
        "00000000",
        -- [0x27] x
        "00000000",
        "00000000",
        "11000110",
        "01101100",
        "00111000",
        "01101100",
        "11000110",
        "00000000",
     	-- [0x28] z
        "00000000",
        "00000000",
        "11111100",
        "10011000",
        "00110000",
        "01100100",
        "11111100",
        "00000000",
     	-- [0x29] space
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
      	-- [0x2A] horizontal border
        "00000000",
        "00000000",
        "00000000",
        "11111111",
        "11111111",
        "00000000",
        "00000000",
        "00000000",
     	-- [0x2B] vertical border
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
    	-- [0x2C] top-left corner
        "00000000",
        "00000000",
        "00000000",
        "00011111",
        "00011111",
        "00011000",
        "00011000",
        "00011000",
    	--- [0x2D] top-right corner
        "00000000",
        "00000000",
        "00000000",
        "11111000",
        "11111000",
        "00011000",
        "00011000",
        "00011000",
    	--- [0x2E] bottom-left corner
        "00011000",
        "00011000",
        "00011000",
        "00011111",
        "00011111",
        "00000000",
        "00000000",
        "00000000",
    	--- [0x2F] bottom-right corner
        "00011000",
        "00011000",
        "00011000",
        "11111000",
        "11111000",
        "00000000",
        "00000000",
        "00000000"
    );
                
begin

    data_o <= rom(to_integer(unsigned(row_i)));

end behavioral;
