library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

use work.constants.all;

entity load_store_unit is
	generic (ADDRESS_WIDTH : NATURAL := 14);
	port (
		clk_i : in STD_LOGIC;
		rst_i : in STD_LOGIC;
		exception_i : in STD_LOGIC;
		mem_req_i : in MEMORY_REQUEST;
		MAR_i : in STD_LOGIC_VECTOR (ADDRESS_WIDTH - 1 downto 0);
		cache_req_o : out CACHE_REQUEST (MAR(ADDRESS_WIDTH - 1 downto 0));
		unaligned_access_o : out STD_LOGIC;
		data_i : in STD_LOGIC_VECTOR (63 downto 0);
		data_o : out STD_LOGIC_VECTOR (63 downto 0));
end load_store_unit;

architecture behavioral of load_store_unit is

	signal we : STD_LOGIC_VECTOR (7 downto 0);
	signal unaligned_access, unaligned, is_signed : STD_LOGIC := '0';
	signal reg_data, data_mem : STD_LOGIC_VECTOR (63 downto 0);

	signal b : STD_LOGIC_VECTOR (7 downto 0);
	signal h : STD_LOGIC_VECTOR (15 downto 0);
	signal w : STD_LOGIC_VECTOR (31 downto 0);
	signal lb, lh, lw, d, MDR : STD_LOGIC_VECTOR (63 downto 0);
	signal unaligned_address, unaligned_address_reg : STD_LOGIC_VECTOR (ADDRESS_WIDTH - 1 downto 0);
    signal halfword_unaligned : STD_LOGIC;
    signal int_column : integer range 0 to 7;
    
    alias column : STD_LOGIC_VECTOR (2 downto 0) is MAR_i(2 downto 0);
    
begin

	CHECK_UNALIGNED : process (mem_req_i.MEMOp, MAR_i)
	begin
		unaligned <= '0';
		case mem_req_i.MEMOp is
			when LSU_LH | LSU_LHU | LSU_SH => unaligned <= and column;
			when LSU_LW | LSU_LWU | LSU_SW => unaligned <= column(2) and (or column(1 downto 0));
			when LSU_LD | LSU_SD => unaligned <= or column;
			when others => unaligned <= '0';
		end case;
	end process;

    int_column <= to_integer(unsigned(MAR_i(2 downto 0)));
	BYTE_SELECT : process (all)
	begin
	    we <= (others => '0');
        case mem_req_i.MEMOp is
            when LSU_SB => we(int_column) <= '1';
            when LSU_SH =>
                if unaligned_access = '0' then
                    we(int_column + 1 downto int_column) <= "11";
                else
                    we <= X"01";
                end if;
            when LSU_SW =>
                if unaligned_access = '0' then
                    we(int_column + 3 downto int_column) <= "1111";
                else
                    case int_column is
                        when 5 => we <= X"01";
                        when 6 => we <= X"03";
                        when others => we <= X"07";
                    end case;
                end if;
            when LSU_SD =>
                if unaligned_access = '0' then
                    we <= (others => '1');
                else
                    case int_column is
                        when 1 => we <= X"01";
                        when 2 => we <= X"03";
                        when 3 => we <= X"07";
                        when 4 => we <= X"0F";
                        when 5 => we <= X"1F";
                        when 6 => we <= X"3F";
                        when 7 => we <= X"7F";
                        when others => we <= X"00";
                    end case;
                end if;
            when others => we <= X"00";
        end case;
	end process;

	MDR_SELECT : process (column, mem_req_i.MDR)
	begin
		case column is
			when "000" => MDR <= mem_req_i.MDR;
			when "001" => MDR <= mem_req_i.MDR(55 downto 0) & mem_req_i.MDR(63 downto 56);
			when "010" => MDR <= mem_req_i.MDR(47 downto 0) & mem_req_i.MDR(63 downto 48);
			when "011" => MDR <= mem_req_i.MDR(39 downto 0) & mem_req_i.MDR(63 downto 40);
			when "100" => MDR <= mem_req_i.MDR(31 downto 0) & mem_req_i.MDR(63 downto 32);
			when "101" => MDR <= mem_req_i.MDR(23 downto 0) & mem_req_i.MDR(63 downto 24);
			when "110" => MDR <= mem_req_i.MDR(15 downto 0) & mem_req_i.MDR(63 downto 16);
			when "111" => MDR <= mem_req_i.MDR(7 downto 0) & mem_req_i.MDR(63 downto 8);
			when others => MDR <= (others => '0'); 
		end case;
	end process;

	DATA_REGISTER : process (clk_i)
	begin
		if rising_edge(clk_i) then
			if unaligned = '1' then
				reg_data <= data_i;
			end if;
		end if;
	end process;

	process (clk_i)
	begin
		if rising_edge(clk_i) then
			if rst_i = '1' or exception_i = '1' then
				unaligned_access <= '0';
			else
			     if unaligned_access = '1' then
			        unaligned_access <= '0';
			     elsif unaligned = '1' then
                    unaligned_access <= '1';
                    unaligned_address_reg <= unaligned_address;
                 end if;
			end if;
		end if;
	end process;
 	
    with column select
        b <= data_i(7 downto 0) when "000",
             data_i(15 downto 8) when "001",
             data_i(23 downto 16) when "010",
             data_i(31 downto 24) when "011",
             data_i(39 downto 32) when "100",
             data_i(47 downto 40) when "101",
             data_i(55 downto 48) when "110",
	         data_i(63 downto 56) when "111",
	         (others => '0') when others;	    	

    with column select
        h <= data_i(15 downto 0) when "000",
             data_i(23 downto 8) when "001",
             data_i(31 downto 16) when "010",
             data_i(39 downto 24) when "011",
             data_i(47 downto 32) when "100",
             data_i(55 downto 40) when "101",
             data_i(63 downto 48) when "110",
             data_i(7 downto 0) & reg_data(63 downto 56) when "111",
	         (others => '0') when others;	
	  

	with column select 
        w <= data_i(31 downto 0) when "000",
             data_i(39 downto 8) when "001",
             data_i(47 downto 16) when "010",
             data_i(55 downto 24) when "011",
             data_i(63 downto 32) when "100",
--             data(71 downto 40) when "101",
--             data(79 downto 48) when "110",
--             data(87 downto 56) when "111",
             (others => '0') when others;
	
    with column select 
        d <= data_i when "000",
--             data(71 downto 8) when "001",
--             data(79 downto 16) when "010",
--             data(87 downto 24) when "011",
--             data(95 downto 32) when "100",
--             data(103 downto 40) when "101",
--             data(111 downto 48) when "110",
--             data(119 downto 56) when "111",
             (others => '0') when others;
             
	with mem_req_i.MEMOp select
	   is_signed <= '1' when LSU_LB | LSU_LH | LSU_LW,
	 	            '0' when others;
	
    lb <= (63 downto 8 => ( b(7) and is_signed ) ) & b;
	lh <= (63 downto 16 => ( h(15) and is_signed ) ) & h;
	lw <= (63 downto 32 => ( w(31) and is_signed ) ) & w;

	with mem_req_i.MEMOp select
	   data_mem <= lb when LSU_LB | LSU_LBU,
		           lh when LSU_LH | LSU_LHU,
		           lw when LSU_LW | LSU_LWU,
		           d when LSU_LD,
		           (others => '0') when others;


    unaligned_address <= STD_LOGIC_VECTOR(unsigned(MAR_i) + 1);
	unaligned_access_o <= unaligned and (not unaligned_access);
	
	data_o <= data_mem when mem_req_i.enable_mem else (others => '0');
	
	cache_req_o.MAR <= MAR_i when unaligned_access = '0' else unaligned_address_reg;

	cache_req_o.MDR <= MDR;
	cache_req_o.we <= we;

end behavioral;